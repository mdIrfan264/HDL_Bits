module top_module( input in, output out );

  // just assign the output with the negation of input
    assign out = ~in;
endmodule
