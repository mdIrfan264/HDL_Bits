module top_module( input in, output out );

  // assign the output variable with the input
   assign out = in;

endmodule
