module top_module(
    output zero
);
  // Module body starts after semicolon
  // just assign output variable low
  
assign zero = 1'b0;
endmodule
