module top_module( output one );

// Insert your code here
//just assign output variable high
    assign one = 1'b1;

endmodule
