module top_module( 
    input a, 
    input b, 
    output out );
  //just assign the output with AND gate operation of two input
    assign out = a&b;

endmodule
